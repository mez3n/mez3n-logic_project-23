module sbox (output reg [7:0] out,input [7:0] in);

  always @* begin
    case (in)
8'h	00	: out = 8'h	63	;
8'h	01	: out = 8'h	7C	;
8'h	02	: out = 8'h	77	;
8'h	03	: out = 8'h	7B	;
8'h	04	: out = 8'h	F2	;
8'h	05	: out = 8'h	6B	;
8'h	06	: out = 8'h	6F	;
8'h	07	: out = 8'h	C5	;
8'h	08	: out = 8'h	30	;
8'h	09	: out = 8'h	01	;
8'h	0A	: out = 8'h	67	;
8'h	0B	: out = 8'h	2B	;
8'h	0C	: out = 8'h	FE	;
8'h	0D	: out = 8'h	D7	;
8'h	0E	: out = 8'h	AB	;
8'h	0F	: out = 8'h	76	;
8'h	10	: out = 8'h	CA	;
8'h	11	: out = 8'h	82	;
8'h	12	: out = 8'h	C9	;
8'h	13	: out = 8'h	7D	;
8'h	14	: out = 8'h	FA	;
8'h	15	: out = 8'h	59	;
8'h	16	: out = 8'h	47	;
8'h	17	: out = 8'h	F0	;
8'h	18	: out = 8'h	AD	;
8'h	19	: out = 8'h	D4	;
8'h	1A	: out = 8'h	A2	;
8'h	1B	: out = 8'h	AF	;
8'h	1C	: out = 8'h	9C	;
8'h	1D	: out = 8'h	A4	;
8'h	1E	: out = 8'h	72	;
8'h	1F	: out = 8'h	C0	;
8'h	20	: out = 8'h	B7	;
8'h	21	: out = 8'h	FD	;
8'h	22	: out = 8'h	93	;
8'h	23	: out = 8'h	26	;
8'h	24	: out = 8'h	36	;
8'h	25	: out = 8'h	3F	;
8'h	26	: out = 8'h	F7	;
8'h	27	: out = 8'h	CC	;
8'h	28	: out = 8'h	34	;
8'h	29	: out = 8'h	A5	;
8'h	2A	: out = 8'h	E5	;
8'h	2B	: out = 8'h	F1	;
8'h	2C	: out = 8'h	71	;
8'h	2D	: out = 8'h	D8	;
8'h	2E	: out = 8'h	31	;
8'h	2F	: out = 8'h	15	;
8'h	30	: out = 8'h	04	;
8'h	31	: out = 8'h	C7	;
8'h	32	: out = 8'h	23	;
8'h	33	: out = 8'h	C3	;
8'h	34	: out = 8'h	18	;
8'h	35	: out = 8'h	96	;
8'h	36	: out = 8'h	05	;
8'h	37	: out = 8'h	9A	;
8'h	38	: out = 8'h	07	;
8'h	39	: out = 8'h	12	;
8'h	3A	: out = 8'h	80	;
8'h	3B	: out = 8'h	E2	;
8'h	3C	: out = 8'h	EB	;
8'h	3D	: out = 8'h	27	;
8'h	3E	: out = 8'h	B2	;
8'h	3F	: out = 8'h	75	;
8'h	40	: out = 8'h	09	;
8'h	41	: out = 8'h	83	;
8'h	42	: out = 8'h	2C	;
8'h	43	: out = 8'h	1A	;
8'h	44	: out = 8'h	1B	;
8'h	45	: out = 8'h	6E	;
8'h	46	: out = 8'h	5A	;
8'h	47	: out = 8'h	A0	;
8'h	48	: out = 8'h	52	;
8'h	49	: out = 8'h	3B	;
8'h	4A	: out = 8'h	D6	;
8'h	4B	: out = 8'h	B3	;
8'h	4C	: out = 8'h	29	;
8'h	4D	: out = 8'h	E3	;
8'h	4E	: out = 8'h	2F	;
8'h	4F	: out = 8'h	84	;
8'h	50	: out = 8'h	53	;
8'h	51	: out = 8'h	D1	;
8'h	52	: out = 8'h	00	;
8'h	53	: out = 8'h	ED	;
8'h	54	: out = 8'h	20	;
8'h	55	: out = 8'h	FC	;
8'h	56	: out = 8'h	B1	;
8'h	57	: out = 8'h	5B	;
8'h	58	: out = 8'h	6A	;
8'h	59	: out = 8'h	CB	;
8'h	5A	: out = 8'h	BE	;
8'h	5B	: out = 8'h	39	;
8'h	5C	: out = 8'h	4A	;
8'h	5D	: out = 8'h	4C	;
8'h	5E	: out = 8'h	58	;
8'h	5F	: out = 8'h	CF	;
8'h	60	: out = 8'h	D0	;
8'h	61	: out = 8'h	EF	;
8'h	62	: out = 8'h	AA	;
8'h	63	: out = 8'h	FB	;
8'h	64	: out = 8'h	43	;
8'h	65	: out = 8'h	4D	;
8'h	66	: out = 8'h	33	;
8'h	67	: out = 8'h	85	;
8'h	68	: out = 8'h	45	;
8'h	69	: out = 8'h	F9	;
8'h	6A	: out = 8'h	02	;
8'h	6B	: out = 8'h	7F	;
8'h	6C	: out = 8'h	50	;
8'h	6D	: out = 8'h	3C	;
8'h	6E	: out = 8'h	9F	;
8'h	6F	: out = 8'h	A8	;
8'h	70	: out = 8'h	51	;
8'h	71	: out = 8'h	A3	;
8'h	72	: out = 8'h	40	;
8'h	73	: out = 8'h	8F	;
8'h	74	: out = 8'h	92	;
8'h	75	: out = 8'h	9D	;
8'h	76	: out = 8'h	38	;
8'h	77	: out = 8'h	F5	;
8'h	78	: out = 8'h	BC	;
8'h	79	: out = 8'h	B6	;
8'h	7A	: out = 8'h	DA	;
8'h	7B	: out = 8'h	21	;
8'h	7C	: out = 8'h	10	;
8'h	7D	: out = 8'h	FF	;
8'h	7E	: out = 8'h	F3	;
8'h	7F	: out = 8'h	D2	;
8'h	80	: out = 8'h	CD	;
8'h	81	: out = 8'h	0C	;
8'h	82	: out = 8'h	13	;
8'h	83	: out = 8'h	EC	;
8'h	84	: out = 8'h	5F	;
8'h	85	: out = 8'h	97	;
8'h	86	: out = 8'h	44	;
8'h	87	: out = 8'h	17	;
8'h	88	: out = 8'h	C4	;
8'h	89	: out = 8'h	A7	;
8'h	8A	: out = 8'h	7E	;
8'h	8B	: out = 8'h	3D	;
8'h	8C	: out = 8'h	64	;
8'h	8D	: out = 8'h	5D	;
8'h	8E	: out = 8'h	19	;
8'h	8F	: out = 8'h	73	;
8'h	90	: out = 8'h	60	;
8'h	91	: out = 8'h	81	;
8'h	92	: out = 8'h	4F	;
8'h	93	: out = 8'h	DC	;
8'h	94	: out = 8'h	22	;
8'h	95	: out = 8'h	2A	;
8'h	96	: out = 8'h	90	;
8'h	97	: out = 8'h	88	;
8'h	98	: out = 8'h	46	;
8'h	99	: out = 8'h	EE	;
8'h	9A	: out = 8'h	B8	;
8'h	9B	: out = 8'h	14	;
8'h	9C	: out = 8'h	DE	;
8'h	9D	: out = 8'h	5E	;
8'h	9E	: out = 8'h	0B	;
8'h	9F	: out = 8'h	DB	;
8'h	A0	: out = 8'h	E0	;
8'h	A1	: out = 8'h	32	;
8'h	A2	: out = 8'h	3A	;
8'h	A3	: out = 8'h	0A	;
8'h	A4	: out = 8'h	49	;
8'h	A5	: out = 8'h	06	;
8'h	A6	: out = 8'h	24	;
8'h	A7	: out = 8'h	5C	;
8'h	A8	: out = 8'h	C2	;
8'h	A9	: out = 8'h	D3	;
8'h	AA	: out = 8'h	AC	;
8'h	AB	: out = 8'h	62	;
8'h	AC	: out = 8'h	91	;
8'h	AD	: out = 8'h	95	;
8'h	AE	: out = 8'h	E4	;
8'h	AF	: out = 8'h	79	;
8'h	B0	: out = 8'h	E7	;
8'h	B1	: out = 8'h	C8	;
8'h	B2	: out = 8'h	37	;
8'h	B3	: out = 8'h	6D	;
8'h	B4	: out = 8'h	8D	;
8'h	B5	: out = 8'h	D5	;
8'h	B6	: out = 8'h	4E	;
8'h	B7	: out = 8'h	A9	;
8'h	B8	: out = 8'h	6C	;
8'h	B9	: out = 8'h	56	;
8'h	BA	: out = 8'h	F4	;
8'h	BB	: out = 8'h	EA	;
8'h	BC	: out = 8'h	65	;
8'h	BD	: out = 8'h	7A	;
8'h	BE	: out = 8'h	AE	;
8'h	BF	: out = 8'h	08	;
8'h	C0	: out = 8'h	BA	;
8'h	C1	: out = 8'h	78	;
8'h	C2	: out = 8'h	25	;
8'h	C3	: out = 8'h	2E	;
8'h	C4	: out = 8'h	1C	;
8'h	C5	: out = 8'h	A6	;
8'h	C6	: out = 8'h	B4	;
8'h	C7	: out = 8'h	C6	;
8'h	C8	: out = 8'h	E8	;
8'h	C9	: out = 8'h	DD	;
8'h	CA	: out = 8'h	74	;
8'h	CB	: out = 8'h	1F	;
8'h	CC	: out = 8'h	4B	;
8'h	CD	: out = 8'h	BD	;
8'h	CE	: out = 8'h	8B	;
8'h	CF	: out = 8'h	8A	;
8'h	D0	: out = 8'h	70	;
8'h	D1	: out = 8'h	3E	;
8'h	D2	: out = 8'h	B5	;
8'h	D3	: out = 8'h	66	;
8'h	D4	: out = 8'h	48	;
8'h	D5	: out = 8'h	03	;
8'h	D6	: out = 8'h	F6	;
8'h	D7	: out = 8'h	0E	;
8'h	D8	: out = 8'h	61	;
8'h	D9	: out = 8'h	35	;
8'h	DA	: out = 8'h	57	;
8'h	DB	: out = 8'h	B9	;
8'h	DC	: out = 8'h	86	;
8'h	DD	: out = 8'h	C1	;
8'h	DE	: out = 8'h	1D	;
8'h	DF	: out = 8'h	9E	;
8'h	E0	: out = 8'h	E1	;
8'h	E1	: out = 8'h	F8	;
8'h	E2	: out = 8'h	98	;
8'h	E3	: out = 8'h	11	;
8'h	E4	: out = 8'h	69	;
8'h	E5	: out = 8'h	D9	;
8'h	E6	: out = 8'h	8E	;
8'h	E7	: out = 8'h	94	;
8'h	E8	: out = 8'h	9B	;
8'h	E9	: out = 8'h	1E	;
8'h	EA	: out = 8'h	87	;
8'h	EB	: out = 8'h	E9	;
8'h	EC	: out = 8'h	CE	;
8'h	ED	: out = 8'h	55	;
8'h	EE	: out = 8'h	28	;
8'h	EF	: out = 8'h	DF	;
8'h	F0	: out = 8'h	8C	;
8'h	F1	: out = 8'h	A1	;
8'h	F2	: out = 8'h	89	;
8'h	F3	: out = 8'h	0D	;
8'h	F4	: out = 8'h	BF	;
8'h	F5	: out = 8'h	E6	;
8'h	F6	: out = 8'h	42	;
8'h	F7	: out = 8'h	68	;
8'h	F8	: out = 8'h	41	;
8'h	F9	: out = 8'h	99	;
8'h	FA	: out = 8'h	2D	;
8'h	FB	: out = 8'h	0F	;
8'h	FC	: out = 8'h	B0	;
8'h	FD	: out = 8'h	54	;
8'h	FE	: out = 8'h	BB	;
8'h	FF	: out = 8'h	16	;

      default: out = 8'h00;
    endcase
  end

endmodule
